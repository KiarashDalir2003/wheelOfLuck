library verilog;
use verilog.vl_types.all;
entity CounterTB is
end CounterTB;
