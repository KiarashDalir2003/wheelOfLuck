library verilog;
use verilog.vl_types.all;
entity CounterTestbench is
end CounterTestbench;
